//UART wrapper with register bank and mapping logic 

module uart_ip(
    input clk,
    input rst,

    //AXI INTERFACE 

);

//REGISTER BANK 

//MAPPING LOGIC 


//INSTANTIATION

endmodule 